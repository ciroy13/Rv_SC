module top(

);

endmodule : top